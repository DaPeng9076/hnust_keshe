library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity huowushu is
port(hw1,hw2,hw3,hw4,hw5,hw6:out std_logic_vector(3 downto 0));
end huowushu;

architecture hw of huowushu is

begin
	hw1<="1001";
	hw2<="1001";
	hw3<="1001";
	hw4<="1001";
	hw5<="1001";
	hw6<="1001";

	
end hw;